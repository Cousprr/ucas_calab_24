module mycpu_top(
    input  wire        aclk,
    input  wire        aresetn,
    // read requeset
    // master->slave
    output [ 3:0]   arid,
    output [31:0]   araddr,
    output [ 7:0]   arlen,
    output [ 2:0]   arsize,
    output [ 1:0]   arburst,
    output [ 1:0]   arlock,
    output [ 3:0]   arcache,
    output [ 2:0]   arprot,
    output          arvalid,
    // slave->master
    input           arready,
    // read response
    // slave->master
    input  [ 3:0]   rid,
    input  [31:0]   rdata,
    input  [ 1:0]   rresp,
    input           rlast,
    input           rvalid,
    // master->slave
    output          rready,
    // write request
    // master->slave
    output [ 3:0]   awid,
    output [31:0]   awaddr,
    output [ 7:0]   awlen,
    output [ 2:0]   awsize,
    output [ 1:0]   awburst,
    output [ 1:0]   awlock,
    output [ 3:0]   awcache,
    output [ 2:0]   awprot,
    output          awvalid,
    // slave->master
    input           awready,
    // write data
    // master->slave
    output  [ 3:0]  wid,
    output  [31:0]  wdata,
    output  [ 3:0]  wstrb,
    output          wlast,
    output          wvalid,
    // slave->master
    input           wready,
    // write response
    // slave->master
    input  [ 3:0]   bid,
    input  [ 1:0]   bresp,
    input           bvalid,
    // master->slave
    output          bready,

    // trace debug interface
    output wire [31:0] debug_wb_pc,
    output wire [ 3:0] debug_wb_rf_we,
    output wire [ 4:0] debug_wb_rf_wnum,
    output wire [31:0] debug_wb_rf_wdata
);



    wire ID_allow_in;
    wire IF_to_ID_valid;
    wire [69:0] IF_to_ID_bus;//70
    wire [33:0] ID_to_IF_bus;//34
    wire EXE_allow_in;
    wire ID_to_EXE_valid;
    wire [351:0] ID_to_EXE_bus;
    wire [37:0] WB_to_ID_bus;
    wire EXE_to_MEM_valid;
    wire MEM_allow_in;
    wire [200:0]EXE_to_MEM_bus;
    wire MEM_to_WB_valid;
    wire WB_allow_in;
    //wire MEM_to_WB_bus;
    wire [197:0] MEM_to_WB_bus;
    wire [38:0]EXE_wr_bus;
    wire [38:0]MEM_wr_bus;
    wire csr_we;             //дʹ��
    wire [13:0] csr_num;     //�Ĵ�����(д)
    wire [31:0] csr_wmask;    //д����
    wire [31:0] csr_wvalue;   //д����
    wire [13:0] csr_raddr;    //����ַ
    wire [31:0] csr_rvalue;  //������
    wire [31:0] ex_entry;    //�жϳ�����ڵ�ַ
    wire [31:0] ex_exit;     //�жϳ����˳���ַ
    wire ertn_flush;          //ertnָ��ִ�е���Ч�ź�
    wire has_int;            //�ж���Ч�ź�
    wire wb_ex;               //�쳣�������ź�
    wire [5:0] wb_ecode;
    wire [8:0] wb_esubcode;
    wire [31:0] WB_pc;
    wire MEM_ex;
    wire MEM_ertn;
    wire [16:0] MEM_to_csr_bus;
    wire [16:0] EXE_to_csr_bus;
    wire [16:0] WB_to_csr_bus;
    wire [31:0] wb_badvaddr;
    wire csr_has_int;
    wire ldst_cancel;
    wire            inst_sram_req;
    wire            inst_sram_wr;
    wire  [ 1:0]    inst_sram_size;
    wire  [31:0]    inst_sram_addr;
    wire  [ 3:0]    inst_sram_wstrb;
    wire  [31:0]    inst_sram_wdata;
    wire            inst_sram_addr_ok;
    wire            inst_sram_data_ok;
    wire [31:0]     inst_sram_rdata;
    wire            data_sram_req;
    wire            data_sram_wr;
    wire  [ 1:0]    data_sram_size;
    wire  [31:0]    data_sram_addr;
    wire  [ 3:0]    data_sram_wstrb;
    wire  [31:0]    data_sram_wdata;
    wire            data_sram_addr_ok;
    wire            data_sram_data_ok;
    wire [31:0]     data_sram_rdata;

    wire       tlbrd_we;
    wire       tlbsrch_we;
    wire       tlb_hit;
    wire [ 3:0]tlb_hit_index;
    wire [ 3:0]csr_tlbidx_index;
    wire [18:0]csr_tlbidx_vppn;
    wire [18:0]s0_vppn;
    wire       s0_va_bit12;
    wire [ 9:0]s0_asid;
    wire       s0_found;
    wire [ 3:0]s0_index;
    wire [19:0]s0_ppn;
    wire [ 5:0]s0_ps;
    wire [ 1:0]s0_plv;
    wire [ 1:0]s0_mat;
    wire       s0_d;
    wire       s0_v;
    wire [18:0]s1_vppn;
    wire       s1_va_bit12;
    wire [ 9:0]s1_asid;
    wire       s1_found;
    wire [ 3:0]s1_index;
    wire [19:0]s1_ppn;
    wire [ 5:0]s1_ps;
    wire [ 1:0]s1_plv;
    wire [ 1:0]s1_mat;
    wire       s1_d;
    wire       s1_v;
    wire [ 4:0]invtlb_op;
    wire       invtlb_valid;
    wire       we;
    wire [ 3:0]w_index;
    wire       w_e;
    wire [18:0]w_vppn;
    wire [ 5:0]w_ps;
    wire [ 9:0]w_asid;
    wire       w_g;
    wire [19:0]w_ppn0;
    wire [ 1:0]w_plv0;
    wire [ 1:0]w_mat0;
    wire       w_d0;
    wire       w_v0;
    wire [19:0]w_ppn1;
    wire [ 1:0]w_plv1;
    wire [ 1:0]w_mat1;
    wire       w_d1;
    wire       w_v1;
    wire [ 3:0]r_index;
    wire       r_e;
    wire [18:0]r_vppn;
    wire [ 5:0]r_ps;
    wire [ 9:0]r_asid;
    wire       r_g;
    wire [19:0]r_ppn0;
    wire [ 1:0]r_plv0;
    wire [ 1:0]r_mat0;
    wire       r_d0;
    wire       r_v0;
    wire [19:0]r_ppn1;
    wire [ 1:0]r_plv1;
    wire [ 1:0]r_mat1;
    wire       r_d1;
    wire       r_v1;
    wire [18:0]csr_tlbehi_vppn;
    wire [ 9:0]csr_asid_asid;
    assign s0_asid = csr_asid_asid;

bridge my_bridge(
        .aclk               (aclk      ),
        .aresetn            (aresetn   ),

        .arid               (arid      ),
        .araddr             (araddr    ),
        .arlen              (arlen     ),
        .arsize             (arsize    ),
        .arburst            (arburst   ),
        .arlock             (arlock    ),
        .arcache            (arcache   ),
        .arprot             (arprot    ),
        .arvalid            (arvalid   ),
        .arready            (arready   ),
                    
        .rid                (rid       ),
        .rdata              (rdata     ),
        .rresp              (rresp     ),
        .rlast              (rlast     ),
        .rvalid             (rvalid    ),
        .rready             (rready    ),
                
        .awid               (awid      ),
        .awaddr             (awaddr    ),
        .awlen              (awlen     ),
        .awsize             (awsize    ),
        .awburst            (awburst   ),
        .awlock             (awlock    ),
        .awcache            (awcache   ),
        .awprot             (awprot    ),
        .awvalid            (awvalid   ),
        .awready            (awready   ),
        
        .wid                (wid       ),
        .wdata              (wdata     ),
        .wstrb              (wstrb     ),
        .wlast              (wlast     ),
        .wvalid             (wvalid    ),
        .wready             (wready    ),
        
        .bid                (bid       ),
        .bresp              (bresp     ),
        .bvalid             (bvalid    ),
        .bready             (bready    ),
        .inst_sram_req      (inst_sram_req    ),
        .inst_sram_wr       (inst_sram_wr     ),
        .inst_sram_size     (inst_sram_size   ),
        .inst_sram_wstrb    (inst_sram_wstrb  ),
        .inst_sram_addr     (inst_sram_addr   ),
        .inst_sram_wdata    (inst_sram_wdata  ),
        .inst_sram_addr_ok  (inst_sram_addr_ok),
        .inst_sram_data_ok  (inst_sram_data_ok),
        .inst_sram_rdata    (inst_sram_rdata  ),
        .data_sram_req      (data_sram_req    ),
        .data_sram_wr       (data_sram_wr     ),
        .data_sram_size     (data_sram_size   ),
        .data_sram_addr     (data_sram_addr   ),
        .data_sram_wstrb    (data_sram_wstrb  ),
        .data_sram_wdata    (data_sram_wdata  ),
        .data_sram_addr_ok  (data_sram_addr_ok),
        .data_sram_data_ok  (data_sram_data_ok),
        .data_sram_rdata    (data_sram_rdata  )
    );


    IF u_IF(
    .clk(aclk),
    .resetn(aresetn),
    .ID_allow_in(ID_allow_in),
    .IF_to_ID_valid(IF_to_ID_valid),
    .IF_to_ID_bus(IF_to_ID_bus),//pc & instruction
    .ID_to_IF_bus(ID_to_IF_bus),//br_takan & br_target
    .inst_sram_req(inst_sram_req),
    .inst_sram_wr(inst_sram_wr),
    .inst_sram_size(inst_sram_size),
    .inst_sram_wstrb(inst_sram_wstrb),
    .inst_sram_addr(inst_sram_addr),
    .inst_sram_wdata(inst_sram_wdata),
    .inst_sram_rdata(inst_sram_rdata),
    .inst_sram_addr_ok(inst_sram_addr_ok),
    .inst_sram_data_ok(inst_sram_data_ok),
    .wb_ex(wb_ex),
    .ertn_flush(ertn_flush),
    .ex_entry(ex_entry),
    .ex_exit(ex_exit)
    );
 
    ID u_ID(
    .clk(aclk),
    .resetn(aresetn),
    .IF_to_ID_valid(IF_to_ID_valid),//IF���������������ȷ���
    .ID_allow_in(ID_allow_in),//ID������������
    .IF_to_ID_bus(IF_to_ID_bus),//pc & instruction
    .ID_to_IF_bus(ID_to_IF_bus),//br_takan & br_target
    .EXE_allow_in(EXE_allow_in),
    .ID_to_EXE_valid(ID_to_EXE_valid),
    .ID_to_EXE_bus(ID_to_EXE_bus),
    .WB_to_ID_bus(WB_to_ID_bus),
    .EXE_wr_bus(EXE_wr_bus),
    .MEM_wr_bus(MEM_wr_bus),
    .csr_rvalue(csr_rvalue),
    .csr_raddr(csr_raddr),
    .EXE_to_csr_bus(EXE_to_csr_bus),
    .MEM_to_csr_bus(MEM_to_csr_bus),
    .WB_to_csr_bus(WB_to_csr_bus),
    .csr_has_int(csr_has_int),
    .wb_ex(wb_ex)
    );
    
    EXE u_EXE(
    .clk(aclk),
    .resetn(aresetn),
    .EXE_allow_in(EXE_allow_in),
    .ID_to_EXE_valid(ID_to_EXE_valid),
    .ID_to_EXE_bus(ID_to_EXE_bus),
    .EXE_to_MEM_valid(EXE_to_MEM_valid),
    .MEM_allow_in(MEM_allow_in),
    .EXE_to_MEM_bus(EXE_to_MEM_bus),
    .data_sram_req(data_sram_req),
    .data_sram_wr(data_sram_wr),
    .data_sram_size(data_sram_size),
    .data_sram_wstrb(data_sram_wstrb),
    .data_sram_addr(data_sram_addr),
    .data_sram_wdata(data_sram_wdata),
    .data_sram_addr_ok(data_sram_addr_ok),
    .EXE_wr_bus(EXE_wr_bus),
    .EXE_to_csr_bus(EXE_to_csr_bus),
    .wb_ex(wb_ex),
    .ertn_flush(ertn_flush),
    .MEM_ex(MEM_ex),
    .MEM_ertn(MEM_ertn),
    .ldst_cancel(ldst_cancel),
    .s1_vppn(s1_vppn),
    .s1_va_bit12(s1_va_bit12),
    .s1_asid(s1_asid),
    .s1_found(s1_found),
    .s1_index(s1_index),
    .s1_ppn(s1_ppn),
    .s1_ps(s1_ps),
    .s1_plv(s1_plv),
    .s1_mat(s1_mat),
    .s1_d(s1_d),
    .s1_v(s1_v),
    .invtlb_valid(invtlb_valid),
    .invtlb_op(invtlb_op),
    .csr_asid_asid(csr_asid_asid),
    .csr_tlbehi_vppn(csr_tlbehi_vppn)
    );
    
    MEM u_MEM(
    .clk(aclk),
    .resetn(aresetn),
    .MEM_allow_in(MEM_allow_in),
    .EXE_to_MEM_valid(EXE_to_MEM_valid),
    .EXE_to_MEM_bus(EXE_to_MEM_bus),
    .MEM_to_WB_valid(MEM_to_WB_valid),
    .WB_allow_in(WB_allow_in),
    .MEM_to_WB_bus(MEM_to_WB_bus),
    .data_sram_rdata(data_sram_rdata),
    .data_sram_data_ok(data_sram_data_ok),
    .MEM_wr_bus(MEM_wr_bus),
    .MEM_ex(MEM_ex),
    .MEM_ertn(MEM_ertn),
    .MEM_to_csr_bus(MEM_to_csr_bus),
    .wb_ex(wb_ex),
    .ertn_flush(ertn_flush),
    .ldst_cancel(ldst_cancel)
    );
    WB u_WB(
    .clk(aclk),
    .resetn(aresetn),
    .WB_allow_in(WB_allow_in),
    .MEM_to_WB_valid(MEM_to_WB_valid),
    .MEM_to_WB_bus(MEM_to_WB_bus),
    .WB_to_ID_bus(WB_to_ID_bus),
    .debug_wb_pc(debug_wb_pc),
    .debug_wb_rf_we(debug_wb_rf_we),
    .debug_wb_rf_wnum(debug_wb_rf_wnum),
    .debug_wb_rf_wdata(debug_wb_rf_wdata),
    .csr_we(csr_we),              //дʹ��
    .csr_num(csr_num),      //�Ĵ�����(д)
    .csr_wmask(csr_wmask),    //д����
    .csr_wvalue(csr_wvalue),   //д����
    .wb_ex(wb_ex),               //�쳣�������ź�
    .wb_ecode(wb_ecode),
    .wb_esubcode(wb_esubcode),
    .WB_pc(WB_pc),
    .ertn_flush(ertn_flush),
    .WB_to_csr_bus(WB_to_csr_bus),
    .wb_badvaddr(wb_badvaddr),
    .refetch(refetch),
    .r_index(r_index),
    .tlbrd_we(tlbrd_we),
    .csr_tlbidx_index(csr_tlbidx_index),
    .tlbwr_we(tlbwr_we),
    .tlbfill_we(tlbfill_we),
    .tlbsrch_we(tlbsrch_we),
    .w_index(w_index),
    .tlb_we(we),//tlbwr_we | tlbfill_we
    .tlb_hit(tlb_hit),
    .tlb_hit_index(tlb_hit_index)
    );
    
    csr u_csr(
    .clk(aclk),
    .resetn(aresetn),
    .csr_we(csr_we),              //дʹ��
    .csr_num(csr_num),      //�Ĵ�����(д)
    .csr_wmask(csr_wmask),    //д����
    .csr_wvalue(csr_wvalue),   //д����
    .csr_raddr(csr_raddr),    //����ַ
    .csr_rvalue(csr_rvalue),  //������
    .ex_entry(ex_entry),    //�жϳ�����ڵ�ַ
    .ex_exit(ex_exit),     //�жϳ����˳���ַ
    .ertn_flush(ertn_flush),          //ertnָ��ִ�е���Ч�ź�
    .csr_has_int(csr_has_int),            //�ж���Ч�ź�
    .wb_ex(wb_ex),               //�쳣�������ź�
    .wb_ecode(wb_ecode),
    .wb_esubcode(wb_esubcode),
    .WB_pc(WB_pc),
    .wb_badvaddr(wb_badvaddr),
    .csr_asid_asid(csr_asid_asid),
    .csr_tlbehi_vppn(csr_tlbehi_vppn),
    .csr_tlbidx_index(csr_tlbidx_index),
    .tlbrd_we(tlbrd_we),
    .tlbsrch_we(tlbsrch_we),
    .tlbsrch_hit(tlb_hit),
    .tlb_hit_index(tlb_hit_index),
    .r_tlb_e(r_e),
    .r_tlb_ps(r_ps),
    .r_tlb_vppn(r_vppn),
    .r_tlb_asid(r_asid),
    .r_tlb_g(r_g),
    .r_tlb_ppn0(r_ppn0),
    .r_tlb_plv0(r_plv0),
    .r_tlb_mat0(r_mat0),
    .r_tlb_d0(r_d0),
    .r_tlb_v0(r_v0),
    .r_tlb_ppn1(r_ppn1),
    .r_tlb_plv1(r_plv1),
    .r_tlb_mat1(r_mat1),
    .r_tlb_d1(r_d1),
    .r_tlb_v1(r_v1),
    .w_tlb_e(w_e),
    .w_tlb_ps(w_ps),
    .w_tlb_vppn(w_vppn),
    .w_tlb_asid(w_asid),
    .w_tlb_g(w_g),
    .w_tlb_ppn0(w_ppn0),
    .w_tlb_plv0(w_plv0),
    .w_tlb_mat0(w_mat0),
    .w_tlb_d0(w_d0),
    .w_tlb_v0(w_v0),
    .w_tlb_ppn1(w_ppn1),
    .w_tlb_plv1(w_plv1),
    .w_tlb_mat1(w_mat1),
    .w_tlb_d1(w_d1),
    .w_tlb_v1(w_v1)
    );

    tlb u_tlb(
        .clk(aclk),
        .s0_vppn(s0_vppn),
        .s0_va_bit12(s0_va_bit12),
        .s0_asid(s0_asid),
        .s0_found(s0_found),
        .s0_index(s0_index),
        .s0_ppn(s0_ppn),
        .s0_ps(s0_ps),
        .s0_plv(s0_plv),
        .s0_mat(s0_mat),
        .s0_d(s0_d),
        .s0_v(s0_v),
        .s1_vppn(s1_vppn),
        .s1_va_bit12(s1_va_bit12),
        .s1_asid(s1_asid),
        .s1_found(s1_found),
        .s1_index(s1_index),
        .s1_ppn(s1_ppn),
        .s1_ps(s1_ps),
        .s1_plv(s1_plv),
        .s1_mat(s1_mat),
        .s1_d(s1_d),
        .s1_v(s1_v),
        .invtlb_valid(invtlb_valid),
        .invtlb_op(invtlb_op),
        .we(we),
        .w_index(w_index),
        .w_e(w_e),
        .w_vppn(w_vppn),
        .w_ps(w_ps),
        .w_asid(w_asid),
        .w_g(w_g),
        .w_ppn0(w_ppn0),
        .w_plv0(w_plv0),
        .w_mat0(w_mat0),
        .w_d0(w_d0),
        .w_v0(w_v0),
        .w_ppn1(w_ppn1),
        .w_plv1(w_plv1),
        .w_mat1(w_mat1),
        .w_d1(w_d1),
        .w_v1(w_v1),
        .r_index(r_index),
        .r_e(r_e),
        .r_vppn(r_vppn),
        .r_ps(r_ps),
        .r_asid(r_asid),
        .r_g(r_g),
        .r_ppn0(r_ppn0),
        .r_plv0(r_plv0),
        .r_mat0(r_mat0),
        .r_d0(r_d0),
        .r_v0(r_v0),
        .r_ppn1(r_ppn1),
        .r_plv1(r_plv1),
        .r_mat1(r_mat1),
        .r_d1(r_d1),
        .r_v1(r_v1)
    );
//wire        load_op;

endmodule
